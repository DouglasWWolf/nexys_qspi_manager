
//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 14-Aug-2024  1.0.0  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 14;
localparam VERSION_MONTH = 8;
localparam VERSION_YEAR  = 2024;

localparam RTL_TYPE      = 81424;
localparam RTL_SUBTYPE   = 0;



/*
    After final falling SCK edge, do we need a delay before releasing CS?

*/